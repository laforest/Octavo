
// Selects between data read from RAM and from I/O ports, if I/O was detected
// earlier.

module Read_Select
#(
)
(
);

 // put a couple of addressed muxes here, addressed with the I/O detect output

endmodule


