
// Assembly code precedes.

        $writememh(INIT_FILE, mem, START_ADDR, END_ADDR);
    end

// "endmodule" follows.

